`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:18:05 05/21/2016 
// Design Name: 
// Module Name:    tb_top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tb_top(
    );

parameter ADD    = 4'b0000;
parameter SUB    = 4'b0001;
parameter SHIFT  = 4'b0010;
parameter CMP    = 4'b0011;
parameter EXOR   = 4'b0100;
parameter BCMP   = 4'b0101;
parameter AND    = 4'b0110;
parameter NAND   = 4'b0111;
parameter OR     = 4'b1000;
parameter NOR    = 4'b1001;



endmodule
